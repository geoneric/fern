netcdf earth {
dimensions:
variables:
// global attributes:
data:
}
