netcdf earth {

dimensions:

variables:
    double gravity;

:Conventions = "COARDS";

data:
    gravity = 9.8;
}
